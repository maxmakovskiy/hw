// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Sat Sep 04 00:43:17 2021"

module strongmore(
	a0,
	b0,
	a1,
	b1,
	a2,
	b2,
	a3,
	b3,
	y
);


input wire	a0;
input wire	b0;
input wire	a1;
input wire	b1;
input wire	a2;
input wire	b2;
input wire	a3;
input wire	b3;
output wire	y;

wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;

assign	SYNTHESIZED_WIRE_64 = 1;



assign	SYNTHESIZED_WIRE_58 = a0 ^ SYNTHESIZED_WIRE_63;

assign	SYNTHESIZED_WIRE_51 = a0 & SYNTHESIZED_WIRE_1 & SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_5 =  ~SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_52 = a0 & SYNTHESIZED_WIRE_63 & SYNTHESIZED_WIRE_5;

assign	SYNTHESIZED_WIRE_8 = a1 & SYNTHESIZED_WIRE_65 & SYNTHESIZED_WIRE_66;

assign	SYNTHESIZED_WIRE_68 = SYNTHESIZED_WIRE_8 | SYNTHESIZED_WIRE_9 | SYNTHESIZED_WIRE_10 | SYNTHESIZED_WIRE_11;

assign	SYNTHESIZED_WIRE_12 =  ~a1;

assign	SYNTHESIZED_WIRE_11 = SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_65 & SYNTHESIZED_WIRE_66;

assign	SYNTHESIZED_WIRE_16 =  ~SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_9 = a1 & SYNTHESIZED_WIRE_16 & SYNTHESIZED_WIRE_66;

assign	SYNTHESIZED_WIRE_22 =  ~SYNTHESIZED_WIRE_66;

assign	SYNTHESIZED_WIRE_50 = a0 & SYNTHESIZED_WIRE_63 & SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_10 = a1 & SYNTHESIZED_WIRE_65 & SYNTHESIZED_WIRE_22;

assign	SYNTHESIZED_WIRE_25 = a2 & SYNTHESIZED_WIRE_67 & SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_41 = SYNTHESIZED_WIRE_25 | SYNTHESIZED_WIRE_26 | SYNTHESIZED_WIRE_27 | SYNTHESIZED_WIRE_28;

assign	SYNTHESIZED_WIRE_29 =  ~a2;

assign	SYNTHESIZED_WIRE_28 = SYNTHESIZED_WIRE_29 & SYNTHESIZED_WIRE_67 & SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_33 =  ~SYNTHESIZED_WIRE_67;

assign	SYNTHESIZED_WIRE_26 = a2 & SYNTHESIZED_WIRE_33 & SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_37 =  ~SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_27 = a2 & SYNTHESIZED_WIRE_67 & SYNTHESIZED_WIRE_37;

assign	SYNTHESIZED_WIRE_42 = a3 ^ SYNTHESIZED_WIRE_38;

assign	y = SYNTHESIZED_WIRE_39 & SYNTHESIZED_WIRE_40;

assign	SYNTHESIZED_WIRE_43 = SYNTHESIZED_WIRE_41 ^ SYNTHESIZED_WIRE_42;

assign	SYNTHESIZED_WIRE_63 =  ~b0;

assign	SYNTHESIZED_WIRE_65 =  ~b1;

assign	SYNTHESIZED_WIRE_67 =  ~b2;

assign	SYNTHESIZED_WIRE_38 =  ~b3;

assign	SYNTHESIZED_WIRE_40 =  ~SYNTHESIZED_WIRE_43;

assign	SYNTHESIZED_WIRE_46 = a1 ^ SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_54 = SYNTHESIZED_WIRE_66 ^ SYNTHESIZED_WIRE_46;

assign	SYNTHESIZED_WIRE_49 = a2 ^ SYNTHESIZED_WIRE_67;

assign	SYNTHESIZED_WIRE_55 = SYNTHESIZED_WIRE_68 ^ SYNTHESIZED_WIRE_49;

assign	SYNTHESIZED_WIRE_66 = SYNTHESIZED_WIRE_50 | SYNTHESIZED_WIRE_51 | SYNTHESIZED_WIRE_52 | SYNTHESIZED_WIRE_53;

assign	SYNTHESIZED_WIRE_39 = SYNTHESIZED_WIRE_54 | SYNTHESIZED_WIRE_55 | SYNTHESIZED_WIRE_56;

assign	SYNTHESIZED_WIRE_59 =  ~a0;


assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_64 ^ SYNTHESIZED_WIRE_58;

assign	SYNTHESIZED_WIRE_53 = SYNTHESIZED_WIRE_59 & SYNTHESIZED_WIRE_63 & SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_1 =  ~SYNTHESIZED_WIRE_63;


endmodule
